`timescale 1 ps / 1 ps

module part1 (CLOCK_50, CLOCK2_50, KEY, SW, FPGA_I2C_SCLK, FPGA_I2C_SDAT, AUD_XCK, 
		        AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK, AUD_ADCDAT, AUD_DACDAT);

	input CLOCK_50, CLOCK2_50;
	input [0:0] KEY;
	input [9:0]SW;
	// I2C Audio/Video config interface
	output FPGA_I2C_SCLK;
	inout FPGA_I2C_SDAT;
	// Audio CODEC
	output AUD_XCK;
	input AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK;
	input AUD_ADCDAT;
	output AUD_DACDAT;
	
	// Local wires.
	wire read_ready, write_ready, read, write;
	wire [23:0] readdata_left, readdata_right;
	wire [23:0] writedata_left, writedata_right;
	wire reset = ~KEY[0];

	/////////////////////////////////
	// Your code goes here 
	/////////////////////////////////
	
	
	/*
	*********************************
	PART 1
	*********************************
	*/
	
//	assign writedata_left = readdata_left;
//	assign writedata_right = readdata_right;
//	assign read = write;
//	assign write = read_ready & write_ready;

	/*
	*********************************
	PART 2
	*********************************
	*/
//	
//	wire [15:0] counterOut;
//	
//	wire [23:0] tone;
//	
//	counter #(.WIDTH(16)) UPCOUNTER(.incr(write), .reset(reset), .clk(CLOCK_50), .out(counterOut));  
//	
//	tonemem TONEMEMORY(.address(counterOut), .clock(CLOCK_50), .data(), .wren(1'b0), .q(tone));
//	
//	
//	assign writedata_left = SW[9] ? tone:readdata_left;
//	assign writedata_right = SW[9] ? tone:readdata_right;
//	assign read = write;
//	assign write = read_ready & write_ready;
	
	/*
	*********************************
	PART 3
	*********************************
	*/
	
	FIR_Filter #(.N(2)) leftFilter(.dataIn(readdata_left), .en(read_ready & write_ready), .reset(reset), .clk(CLOCK_50), .dataOut(writedata_left));
	FIR_Filter #(.N(2)) rightFilter(.dataIn(readdata_right), .en(read_ready & write_ready), .reset(reset), .clk(CLOCK_50), .dataOut(writedata_right));
	assign read = write;
	assign write = read_ready & write_ready;
/////////////////////////////////////////////////////////////////////////////////
// Audio CODEC interface. 
//
// The interface consists of the following wires:
// read_ready, write_ready - CODEC ready for read/write operation 
// readdata_left, readdata_right - left and right channel data from the CODEC
// read - send data from the CODEC (both channels)
// writedata_left, writedata_right - left and right channel data to the CODEC
// write - send data to the CODEC (both channels)
// AUD_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio CODEC
// I2C_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio/Video Config module
/////////////////////////////////////////////////////////////////////////////////
	clock_generator my_clock_gen(
		// inputs
		CLOCK2_50,
		reset,

		// outputs
		AUD_XCK
	);

	audio_and_video_config cfg(
		// Inputs
		CLOCK_50,
		reset,

		// Bidirectionals
		FPGA_I2C_SDAT,
		FPGA_I2C_SCLK
	);

	audio_codec codec(
		// Inputs
		CLOCK_50,
		reset,

		read,	write,
		writedata_left, writedata_right,

		AUD_ADCDAT,

		// Bidirectionals
		AUD_BCLK,
		AUD_ADCLRCK,
		AUD_DACLRCK,

		// Outputs
		read_ready, write_ready,
		readdata_left, readdata_right,
		AUD_DACDAT
	);

endmodule


